module risc_v_tb ();
  
reg                 CLK_tb;
reg                 RST_tb;



initial 
begin
CLK_tb =1'b0;
RST_tb =1'b0;

#3
RST_tb = 1'b1;

#500
$stop;
end



////////////////////////////////////////// Clock Generator //////////////////////////////////////
always #5 CLK_tb = ~CLK_tb;
////////////////////////////////////////////////////////////////////////////////////////////////





//////////////////////////////////// port maping for design under test /////////////////////////
risc_v DUT(
.CLK(CLK_tb),
.RST(RST_tb)
);

////////////////////////////////////////////////////////////////////////////////////////////////
endmodule